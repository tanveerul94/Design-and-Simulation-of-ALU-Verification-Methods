`include "transaction.sv"
`include "sequence.sv"

//Define sequencer
typedef uvm_sequencer#(alu_transaction) alu_sequencer;