class transaction;
	rand bit[7:0] a;
	rand bit[7:0] b;
	rand bit[3:0] s;
	bit[15:0] out;

endclass:transaction
